module Instrcution (
    input [15:0]a,
    input [15:0]b,
    input cin,
    output [15:0]sum,
    output carry
    );
    wire [16:0]w0,x0;
    wire [16:0]w1,x1;
    wire [16:0]w2,x2;
    wire [16:0]w3,x3;
    wire [16:0]w4,x4;
    wire [16:0]w5,x5;

    //00
    assign w0[0]= cin;
    assign x0[0]= cin;
    assign w0[1]= a[0]&b[0];
    assign x0[1]= a[0]|b[0];
    assign w0[2]= a[1]&b[1];
    assign x0[2]= a[1]|b[1];
    assign w0[3]= a[2]&b[2];
    assign x0[3]= a[2]|b[2];
    assign w0[4]= a[3]&b[3];
    assign x0[4]= a[3]|b[3];
    assign w0[5]= a[4]&b[4];
    assign x0[5]= a[4]|b[4];
    assign w0[6]= a[5]&b[5];
    assign x0[6]= a[5]|b[5];
    assign w0[7]= a[6]&b[6];
    assign x0[7]= a[6]|b[6];
    assign w0[8]= a[7]&b[7];
    assign x0[8]= a[7]|b[7];
    assign w0[9]= a[8]&b[8];
    assign x0[9]= a[8]|b[8];
    assign w0[10]= a[9]&b[9];
    assign x0[10]= a[9]|b[9];
    assign w0[11]= a[10]&b[10];
    assign x0[11]= a[10]|b[10];
    assign w0[12]= a[11]&b[11];
    assign x0[12]= a[11]|b[11];
    assign w0[13]= a[12]&b[12];
    assign x0[13]= a[12]|b[12];
    assign w0[14]= a[13]&b[13];
    assign x0[14]= a[13]|b[13];
    assign w0[15]= a[14]&b[14];
    assign x0[15]= a[14]|b[14];
    assign w0[16]= a[15]&b[15];
    assign x0[16]= a[15]|b[15];

    //1-1
    //x1=wa+ba;
    //x0=wa+za;
    assign w1[0]= w0[0];
    assign x1[0]= x0[0];
    assign w1[1]= (w0[1]&x0[1]) | (w0[0]&x0[1]);
    assign x1[1]= (w0[1]&x0[1]) | (x0[0]&x0[1]);
    assign w1[2]= (w0[2]&x0[2]) | (w0[1]&x0[2]);
    assign x1[2]= (w0[2]&x0[2]) | (x0[1]&x0[2]);
    assign w1[3]= (w0[3]&x0[3]) | (w0[2]&x0[3]);
    assign x1[3]= (w0[3]&x0[3]) | (x0[2]&x0[3]);
    assign w1[4]= (w0[4]&x0[4]) | (w0[3]&x0[4]);
    assign x1[4]= (w0[4]&x0[4]) | (x0[3]&x0[4]);
    assign w1[5]= (w0[5]&x0[5]) | (w0[4]&x0[5]);
    assign x1[5]= (w0[5]&x0[5]) | (x0[4]&x0[5]);
    assign w1[6]= (w0[6]&x0[6]) | (w0[5]&x0[6]);
    assign x1[6]= (w0[6]&x0[6]) | (x0[5]&x0[6]);
    assign w1[7]= (w0[7]&x0[7]) | (w0[6]&x0[7]);
    assign x1[7]= (w0[7]&x0[7]) | (x0[6]&x0[7]);
    assign w1[8]= (w0[8]&x0[8]) | (w0[7]&x0[8]);
    assign x1[8]= (w0[8]&x0[8]) | (x0[7]&x0[8]);
    assign w1[9]= (w0[9]&x0[9]) | (w0[8]&x0[9]);
    assign x1[9]= (w0[9]&x0[9]) | (x0[8]&x0[9]);
    assign w1[10]= (w0[10]&x0[10]) | (w0[9]&x0[10]);
    assign x1[10]= (w0[10]&x0[10]) | (x0[9]&x0[10]);
    assign w1[11]= (w0[11]&x0[11]) | (w0[10]&x0[11]);
    assign x1[11]= (w0[11]&x0[11]) | (x0[10]&x0[11]);
    assign w1[12]= (w0[12]&x0[12]) | (w0[11]&x0[12]);
    assign x1[12]= (w0[12]&x0[12]) | (x0[11]&x0[12]);
    assign w1[13]= (w0[13]&x0[13]) | (w0[12]&x0[13]);
    assign x1[13]= (w0[13]&x0[13]) | (x0[12]&x0[13]);
    assign w1[14]= (w0[14]&x0[14]) | (w0[13]&x0[14]);
    assign x1[14]= (w0[14]&x0[14]) | (x0[13]&x0[14]);
    assign w1[15]= (w0[15]&x0[15]) | (w0[14]&x0[15]);
    assign x1[15]= (w0[15]&x0[15]) | (x0[14]&x0[15]);
    assign w1[16]= (w0[16]&x0[16]) | (w0[15]&x0[16]);
    assign x1[16]= (w0[16]&x0[16]) | (x0[15]&x0[16]);
    //2-2
    assign w2[0]= w1[0];
    assign x2[0]= x1[0];
    assign w2[1]= w1[1];
    assign x2[1]= x1[1];
    assign w2[2]= (w1[2]&x1[2]) | (w1[0]&x1[2]);
    assign x2[2]= (w1[2]&x1[2]) | (x1[0]&x1[2]);
    assign w2[3]= (w1[3]&x1[3]) | (w1[1]&x1[3]);
    assign x2[3]= (w1[3]&x1[3]) | (x1[1]&x1[3]);
    assign w2[4]= (w1[4]&x1[4]) | (w1[2]&x1[4]);
    assign x2[4]= (w1[4]&x1[4]) | (x1[2]&x1[4]);
    assign w2[5]= (w1[5]&x1[5]) | (w1[3]&x1[5]);
    assign x2[5]= (w1[5]&x1[5]) | (x1[3]&x1[5]);
    assign w2[6]= (w1[6]&x1[6]) | (w1[4]&x1[6]);
    assign x2[6]= (w1[6]&x1[6]) | (x1[4]&x1[6]);
    assign w2[7]= (w1[7]&x1[7]) | (w1[5]&x1[7]);
    assign x2[7]= (w1[7]&x1[7]) | (x1[5]&x1[7]);
    assign w2[8]= (w1[8]&x1[8]) | (w1[6]&x1[8]);
    assign x2[8]= (w1[8]&x1[8]) | (x1[6]&x1[8]);
    assign w2[9]= (w1[9]&x1[9]) | (w1[7]&x1[9]);
    assign x2[9]= (w1[9]&x1[9]) | (x1[7]&x1[9]);
    assign w2[10]= (w1[10]&x1[10]) | (w1[8]&x1[10]);
    assign x2[10]= (w1[10]&x1[10]) | (x1[8]&x1[10]);
    assign w2[11]= (w1[11]&x1[11]) | (w1[9]&x1[11]);
    assign x2[11]= (w1[11]&x1[11]) | (x1[9]&x1[11]);
    assign w2[12]= (w1[12]&x1[12]) | (w1[10]&x1[12]);
    assign x2[12]= (w1[12]&x1[12]) | (x1[10]&x1[12]);
    assign w2[13]= (w1[13]&x1[13]) | (w1[11]&x1[13]);
    assign x2[13]= (w1[13]&x1[13]) | (x1[11]&x1[13]);
    assign w2[14]= (w1[14]&x1[14]) | (w1[12]&x1[14]);
    assign x2[14]= (w1[14]&x1[14]) | (x1[12]&x1[14]);
    assign w2[15]= (w1[15]&x1[15]) | (w1[13]&x1[15]);
    assign x2[15]= (w1[15]&x1[15]) | (x1[13]&x1[15]);
    assign w2[16]= (w1[16]&x1[16]) | (w1[14]&x1[16]);
    assign x2[16]= (w1[16]&x1[16]) | (x1[14]&x1[16]);
    //4-4
    assign w3[0]= w2[0];
    assign x3[0]= x2[0];
    assign w3[1]= w2[1];
    assign x3[1]= x2[1];
    assign w3[2]= w2[2];
    assign x3[2]= x2[2];
    assign w3[3]= w2[3];
    assign x3[3]= x2[3];
    assign w3[4]= (w2[4]&x2[4]) | (w2[0]&x2[4]);
    assign x3[4]= (w2[4]&x2[4]) | (x2[0]&x2[4]);
    assign w3[5]= (w2[5]&x2[5]) | (w2[1]&x2[5]);
    assign x3[5]= (w2[5]&x2[5]) | (x2[1]&x2[5]);
    assign w3[6]= (w2[6]&x2[6]) | (w2[2]&x2[6]);
    assign x3[6]= (w2[6]&x2[6]) | (x2[2]&x2[6]);
    assign w3[7]= (w2[7]&x2[7]) | (w2[3]&x2[7]);
    assign x3[7]= (w2[7]&x2[7]) | (x2[3]&x2[7]);
    assign w3[8]= (w2[8]&x2[8]) | (w2[4]&x2[8]);
    assign x3[8]= (w2[8]&x2[8]) | (x2[4]&x2[8]);
    assign w3[9]= (w2[9]&x2[9]) | (w2[5]&x2[9]);
    assign x3[9]= (w2[9]&x2[9]) | (x2[5]&x2[9]);
    assign w3[10]= (w2[10]&x2[10]) | (w2[8]&x2[10]);
    assign x3[10]= (w2[10]&x2[10]) | (x2[8]&x2[10]);
    assign w3[11]= (w2[11]&x2[11]) | (w2[9]&x2[11]);
    assign x3[11]= (w2[11]&x2[11]) | (x2[9]&x2[11]);
    assign w3[12]= (w2[12]&x2[12]) | (w2[10]&x2[12]);
    assign x3[12]= (w2[12]&x2[12]) | (x2[10]&x2[12]);
    assign w3[13]= (w2[13]&x2[13]) | (w2[11]&x2[13]);
    assign x3[13]= (w2[13]&x2[13]) | (x2[11]&x2[13]);
    assign w3[14]= (w2[14]&x2[14]) | (w2[12]&x2[14]);
    assign x3[14]= (w2[14]&x2[14]) | (x2[12]&x2[14]);
    assign w3[15]= (w2[15]&x2[15]) | (w2[13]&x2[15]);
    assign x3[15]= (w2[15]&x2[15]) | (x2[13]&x2[15]);
    assign w3[16]= (w2[16]&x2[16]) | (w2[14]&x2[16]);
    assign x3[16]= (w2[16]&x2[16]) | (x2[14]&x2[16]);
    //8-8
    assign w4[0]= w3[0];
    assign x4[0]= x3[0];
    assign w4[1]= w3[1];
    assign x4[1]= x3[1];
    assign w4[2]= w3[2];
    assign x4[2]= x3[2];
    assign w4[3]= w3[3];
    assign x4[3]= x3[3];
    assign w4[4]= w3[4];
    assign x4[4]= x3[4];
    assign w4[5]= w3[5];
    assign x4[5]= x3[5];
    assign w4[6]= w3[6];
    assign x4[6]= x3[6];
    assign w4[7]= w3[7];
    assign x4[7]= x3[7];
    assign w4[8]= (w3[8]&x3[8]) | (w3[0]&x3[8]);
    assign x4[8]= (w3[8]&x3[8]) | (x3[0]&x3[8]);
    assign w4[9]= (w3[9]&x3[9]) | (w3[1]&x3[9]);
    assign x4[9]= (w3[9]&x3[9]) | (x3[1]&x3[9]);
    assign w4[10]= (w3[10]&x3[10]) | (w3[2]&x3[10]);
    assign x4[10]= (w3[10]&x3[10]) | (x3[2]&x3[10]);
    assign w4[11]= (w3[11]&x3[11]) | (w3[3]&x3[11]);
    assign x4[11]= (w3[11]&x3[11]) | (x3[3]&x3[11]);
    assign w4[12]= (w3[12]&x3[12]) | (w3[4]&x3[12]);
    assign x4[12]= (w3[12]&x3[12]) | (x3[4]&x3[12]);
    assign w4[13]= (w3[13]&x3[13]) | (w3[5]&x3[13]);
    assign x4[13]= (w3[13]&x3[13]) | (x3[5]&x3[13]);
    assign w4[14]= (w3[14]&x3[14]) | (w3[6]&x3[14]);
    assign x4[14]= (w3[14]&x3[14]) | (x3[6]&x3[14]);
    assign w4[15]= (w3[15]&x3[15]) | (w3[7]&x3[15]);
    assign x4[15]= (w3[15]&x3[15]) | (x3[7]&x3[15]);
    assign w4[16]= (w3[16]&x3[16]) | (w3[8]&x3[16]);
    assign x4[16]= (w3[16]&x3[16]) | (x3[8]&x3[16]);
    //16-16
    assign w5[0]= w4[0];
    assign x5[0]= x4[0];
    assign w5[1]= w4[1];
    assign x5[1]= x4[1];
    assign w5[2]= w4[2];
    assign x5[2]= x4[2];
    assign w5[3]= w4[3];
    assign x5[3]= x4[3];
    assign w5[4]= w4[4];
    assign x5[4]= x4[4];
    assign w5[5]= w4[5];
    assign x5[5]= x4[5];
    assign w5[6]= w4[6];
    assign x5[6]= x4[6];
    assign w5[7]= w4[7];
    assign x5[7]= x4[7];
    assign w5[8]= w4[8];
    assign x5[8]= x4[8];
    assign w5[9]= w4[9];
    assign x5[9]= x4[9];
    assign w5[10]= w4[10];
    assign x5[10]= x4[10];
    assign w5[11]= w4[11];
    assign x5[11]= x4[11];
    assign w5[12]= w4[12];
    assign x5[12]= x4[12];
    assign w5[13]= w4[13];
    assign x5[13]= x4[13];
    assign w5[14]= w4[14];
    assign x5[14]= x4[14];
    assign w5[15]= w4[15];
    assign x5[15]= x4[15];
    assign w5[16]= (w4[16]&x4[16]) | (w4[0]&x4[16]);
    assign x5[16]= (w4[16]&x4[16]) | (x4[0]&x4[16]);



    assign sum[0] = a[0]^b[0]^(w5[0]&x5[0]);
    assign sum[1] = a[1]^b[1]^(w5[1]&x5[1]);
    assign sum[2] = a[2]^b[2]^(w5[2]&x5[2]);
    assign sum[3] = a[3]^b[3]^(w5[3]&x5[3]);
    assign sum[4] = a[4]^b[4]^(w5[4]&x5[4]);
    assign sum[5] = a[5]^b[5]^(w5[5]&x5[5]);
    assign sum[6] = a[6]^b[6]^(w5[6]&x5[6]);
    assign sum[7] = a[7]^b[7]^(w5[7]&x5[7]);
    assign sum[8] = a[8]^b[8]^(w5[8]&x5[8]);
    assign sum[9] = a[9]^b[9]^(w5[9]&x5[9]);
    assign sum[10] = a[10]^b[10]^(w5[10]&x5[10]);
    assign sum[11] = a[11]^b[11]^(w5[11]&x5[11]);
    assign sum[12] = a[12]^b[12]^(w5[12]&x5[12]);
    assign sum[13] = a[13]^b[13]^(w5[13]&x5[13]);
    assign sum[14] = a[14]^b[14]^(w5[14]&x5[14]);
    assign sum[15] = a[15]^b[15]^(w5[15]&x5[15]);
    assign carry = (w5[16]&x5[16]);
   
endmodule

